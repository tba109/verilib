///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Tyler Anderson Fri Feb  8 14:58:05 EST 2019
//
// Test for moving sum
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ns

///////////////////////////////////////////////////////////////////////////////////////////////////
// Test cases
///////////////////////////////////////////////////////////////////////////////////////////////////
`define TEST_CASE_1

module tb;
   
   //////////////////////////////////////////////////////////////////////
   // I/O
   //////////////////////////////////////////////////////////////////////   
   parameter CLK_PERIOD = 10;
   reg clk;
   reg rst;

   // Connections
   /*AUTOWIRE*/
   // Beginning of automatic wires (for undeclared instantiated-module outputs)
   wire [23:0]		sum;			// From UUT_0 of moving_sum.v
   // End of automatics
   /*AUTOREGINPUT*/
   // Beginning of automatic reg inputs (for undeclared instantiated-module inputs)
   reg [15:0]		a;			// To UUT_0 of moving_sum.v
   reg [15:0]		b;			// To UUT_0 of moving_sum.v
   reg [31:0]		init_sum;		// To UUT_0 of moving_sum.v
   reg			init_wr;		// To UUT_0 of moving_sum.v
   reg			wr;			// To UUT_0 of moving_sum.v
   // End of automatics
   
   //////////////////////////////////////////////////////////////////////
   // Clock Driver
   //////////////////////////////////////////////////////////////////////
   always @(clk)
     #(CLK_PERIOD / 2.0) clk <= !clk;
				   
   //////////////////////////////////////////////////////////////////////
   // Simulated interfaces
   //////////////////////////////////////////////////////////////////////   
      
   //////////////////////////////////////////////////////////////////////
   // UUT
   //////////////////////////////////////////////////////////////////////   
   moving_sum UUT_0(/*AUTOINST*/
		    // Outputs
		    .sum		(sum[23:0]),
		    // Inputs
		    .clk		(clk),
		    .wr		(wr),
		    .a		(a[15:0]),
		    .b		(b[15:0]),
		    .init_wr	(init_wr),
		    .init_sum	(init_sum[31:0])); 
   

   //////////////////////////////////////////////////////////////////////
   // Test case
   //////////////////////////////////////////////////////////////////////   
   `ifdef TEST_CASE_1
   initial
     begin
	clk = 1'b0;
	rst = 1'b1;
	a <= 0;
	b <= 0;
	init_sum <= 0;
	init_wr <= 0;
	wr <= 0; 
	// Reset	
	#(20* CLK_PERIOD);
	rst = 0; 
	
	// Logging
	$display("");
	$display("------------------------------------------------------");
	$display("Test Case: TEST_CASE_1");

	init_wr = 1;
	init_sum = 16'h2000;
	#(1 * CLK_PERIOD);

	init_wr <= 0;
	b <= 16'h2001;
	wr <= 1; 
	#(1 * CLK_PERIOD);
	wr <= 0; 
	
	init_wr <= 0;
	a <= 16'h2002; 
	b <= 16'h2001;
	wr <= 1; 
	#(1 * CLK_PERIOD);
	wr <= 0; 

	
     end
   `endif

   //////////////////////////////////////////////////////////////////////
   // Tasks (e.g., writing data, etc.)
   //////////////////////////////////////////////////////////////////////   
   
   
   
endmodule

// Local Variables:
// verilog-library-flags:("-y ../")
// End:
   
