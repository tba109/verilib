//////////////////////////////////////////////////////////////////////////////////////////////////
// Tyler Anderson Mon 11/11/2019_14:01:26.20
//
// tb.v
//
//////////////////////////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ns

//////////////////////////////////////////////////////////////////////////////////////////////////
// Test cases
//////////////////////////////////////////////////////////////////////////////////////////////////
`define TEST_CASE_1

module tb;
   
   //////////////////////////////////////////////////////////////////////
   // I/O
   //////////////////////////////////////////////////////////////////////   
   parameter CLK_PERIOD = 10.0;
   reg clk;
   reg rst;

   // Connections
   // Beginning of automatic wires (for undeclared instantiated-module outputs)
   wire			y;			// From OS_0 of one_shot.v
   wire 		busy; 
   // End of automatics
   reg			trig;			// To OS_0 of one_shot.v
   // End of automatics
   
   //////////////////////////////////////////////////////////////////////
   // Clock Driver
   //////////////////////////////////////////////////////////////////////
   always @(clk)
     #(CLK_PERIOD / 2.0) clk <= !clk;
				   
   //////////////////////////////////////////////////////////////////////
   // Simulated interfaces
   //////////////////////////////////////////////////////////////////////   
      
   //////////////////////////////////////////////////////////////////////
   // UUT
   //////////////////////////////////////////////////////////////////////   
   one_shot #(.P_N_WIDTH(32),.P_IO_WIDTH(1))OS_0
     (
      // Outputs
      .y			(y),
      .busy                     (busy), 
      // Inputs
      .clk			(clk),
      .rst_n			(!rst),
      .trig			(trig),
      .n0			(0),
      .n1			(10),
      .a0			(1'b0),
      .a1			(1'b1)); 
   
   //////////////////////////////////////////////////////////////////////
   // Testbench
   //////////////////////////////////////////////////////////////////////   
   initial
     begin
	// Initializations
	clk = 1'b0;
	rst = 1'b1;
     end

   //////////////////////////////////////////////////////////////////////
   // Test case
   //////////////////////////////////////////////////////////////////////   
   `ifdef TEST_CASE_1
   initial
     begin
	trig = 0;
	
	// Reset	
	#(10 * CLK_PERIOD);
	rst = 1'b0;
	#(20* CLK_PERIOD);

	// Logging
	$display("");
	$display("------------------------------------------------------");
	$display("Test Case: TEST_CASE_1");

	// Stimulate UUT
	@(posedge clk) trig = 1; #1;
	@(posedge clk) trig = 0; #1; 

     end
   `endif

   //////////////////////////////////////////////////////////////////////
   // Tasks (e.g., writing data, etc.)
   //////////////////////////////////////////////////////////////////////   
   
   
   
endmodule

// Local Variables:
// verilog-library-flags:("-y ../")
// End:
   
