///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Tyler Anderson Fri Mar 22 12:15:00 EDT 2019
// tb.v
//
// 
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ns

///////////////////////////////////////////////////////////////////////////////////////////////////
// Test cases
///////////////////////////////////////////////////////////////////////////////////////////////////
`define TEST_CASE_1

module tb;
   
   //////////////////////////////////////////////////////////////////////
   // I/O
   //////////////////////////////////////////////////////////////////////   
   parameter CLK_PERIOD = 10;
   reg clk;
   reg rst;

   // Connections
   /*AUTOWIRE*/
   // Beginning of automatic wires (for undeclared instantiated-module outputs)
   wire			valid;			// From IILC_0 of iter_integer_linear_calc.v
   wire [31:0]		y;			// From IILC_0 of iter_integer_linear_calc.v
   // End of automatics
   /*AUTOREGINPUT*/
   // Beginning of automatic reg inputs (for undeclared instantiated-module inputs)
   reg [31:0]		b;			// To IILC_0 of iter_integer_linear_calc.v
   reg [31:0]		m;			// To IILC_0 of iter_integer_linear_calc.v
   reg [31:0]		x;			// To IILC_0 of iter_integer_linear_calc.v
   // End of automatics
   
   //////////////////////////////////////////////////////////////////////
   // Clock Driver
   //////////////////////////////////////////////////////////////////////
   always @(clk)
     #(CLK_PERIOD / 2.0) clk <= !clk;
				   
   //////////////////////////////////////////////////////////////////////
   // Simulated interfaces
   //////////////////////////////////////////////////////////////////////   
      
   //////////////////////////////////////////////////////////////////////
   // UUT
   //////////////////////////////////////////////////////////////////////   
   iter_integer_linear_calc IILC_0(/*AUTOINST*/
				   // Outputs
				   .y			(y[31:0]),
				   .valid		(valid),
				   // Inputs
				   .clk			(clk),
				   .rst			(rst),
				   .m			(m[31:0]),
				   .x			(x[31:0]),
				   .b			(b[31:0])); 
   
   //////////////////////////////////////////////////////////////////////
   // Testbench
   //////////////////////////////////////////////////////////////////////   
   initial
     begin
	// Initializations
	clk = 1'b0;
	rst = 1'b1;
     end

   //////////////////////////////////////////////////////////////////////
   // Test case
   //////////////////////////////////////////////////////////////////////   
   `ifdef TEST_CASE_1
   initial
     begin
	b = 0;
	m = 0;
	x = 0; 
	// Reset	
	#(10 * CLK_PERIOD);
	rst = 1'b0;
	#(20* CLK_PERIOD);

	// Logging
	$display("");
	$display("------------------------------------------------------");
	$display("Test Case: TEST_CASE_1");

	// Stimulate UUT
	b = 10;
	#(10*CLK_PERIOD);
	x = 16;
	m = 11;

	#(100*CLK_PERIOD);
	x = 12;
	m = 7;
	
     end
   `endif

   //////////////////////////////////////////////////////////////////////
   // Tasks (e.g., writing data, etc.)
   //////////////////////////////////////////////////////////////////////   
   
   
   
endmodule

// Local Variables:
// verilog-library-flags:("-y ../")
// End:
   
